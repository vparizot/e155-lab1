
// Onboard LEDs - defining the behavior of 3 LEDS

module top(
	input logic clk, input logic [3:0] s,
	output logic [2:0] led, logic [6:0] seg
);

// variables
	//logic int_osc;
	logic pulse;
	logic led_state = 0;
	logic [24:0] counter = 0;
	logic LEDVAL = 0;

// LED 0 - XOR
	xor (led[0], s[0], s[1]);

// LED 1 - AND
	and (led[1], s[3], s[2]);

// LED 2 - blinks at 2.4 Hz
// Internal high-speed oscillator

	//HSOSC hf_osc (.CLKHFPU(1'b1), .CLKHFEN(1'b1), .CLKHF(int_osc));
	
// Simple clock divider
	always_ff @(posedge clk)
	begin
		counter <= counter + 1;
		// at hz
		if (counter == 10000000)
		begin
			counter <= 0;
			if (LEDVAL == 0) LEDVAL <= 1 ; // turn on LED if off
			else LEDVAL <= 0; //turn OFF led
		end
	end

		 
// Asssign LED outputs
	assign led[2] = LEDVAL;
	
// call other module
always_comb
	begin
		case (s) 
			4'b0000 : seg = 7'b0100011; //1100010; 
			4'b0001 : seg = 7'b1111001; //b1111001;
			4'b0010 : seg = 7'b0100100; //b0010010;
			4'b0011 : seg = 7'b0110000; //b0000110;
			4'b0100 : seg = 7'b0011001; //b1001100;
			4'b0101 : seg = 7'b0010010; //b0100100;
			4'b0110 : seg = 7'b0000010; //b0100000;
			4'b0111 : seg = 7'b1111000; //b0001111;
			4'b1000 : seg = 7'b0000000; //b0000000;
			4'b1001 : seg = 7'b0011000; //b0001100;
			4'b1010 : seg = 7'b0100000; //b0000010;
			4'b1011 : seg = 7'b0000011; //b1100000;
			4'b1100 : seg = 7'b1000110; //b0110001;
			4'b1101 : seg = 7'b0000011; //b1100010;
			4'b1110 : seg = 7'b0000100; //b0010000;
			4'b1111 : seg = 7'b0001110; //b0111000;
			default: seg = 7'b1111111;
		endcase
	end

endmodule